// 32X32 Multiplier test template
module mult32x32_fast_test;

    logic [31:0] a;        // Input a
    logic [31:0] b;        // Input b
    logic start;           // Start signal
    logic [63:0] product;  // Miltiplication product
    logic valid;           // Operation valid indication

    logic clk;             // Clock
    logic reset;           // Reset

// Put your code here
// ------------------

// End of your code

endmodule
